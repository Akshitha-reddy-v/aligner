///////////////////////////////////////////////////////////////////////////////
// File:        cfs_algn_test_pkg.sv
// Author:      Cristian Florin Slav
// Date:        2023-06-27
// Description: Test package.
///////////////////////////////////////////////////////////////////////////////
`ifndef CFS_ALGN_TEST_PKG_SV
  `define CFS_ALGN_TEST_PKG_SV

  `include "uvm_macros.svh"
  //`include "cfs_algn_pkg.sv"

  package cfs_algn_test_pkg;
    import uvm_pkg::*;
    import cfs_algn_pkg::*;
    import cfs_apb_pkg::*;
    import cfs_md_pkg::*;

    `include "cfs_algn_test_defines.sv"
    `include "cfs_algn_test_base.sv"
    `include "cfs_algn_test_reg_access.sv"
    `include "cfs_algn_test_random.sv"
    `include "cfs_algn_test_random_rx_err.sv"

    `include "algn_test_mid_reset.sv"
    `include "algn_test_legal_rx.sv"
    `include "algn_test_illegal_rx.sv"
    `include "algn_test_rxfifo_full.sv"
    `include "algn_test_reg_access.sv"
    `include "algn_test_apb_back2back.sv"
    `include "algn_test_apb_reset_during_access.sv"
    `include "algn_test_split_directed.sv"
    `include "algn_test_legal_rx_ctrl_directed.sv"


  endpackage

`endif
